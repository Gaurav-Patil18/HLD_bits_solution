// Problem: 44 - exams/m2014_q4h
module top_module (
    input in,
    output out);
assign out=in;
endmodule
