// Problem: 1 - step_one

module top_module( output one );

// Insert your code here
    assign one = 1;

endmodule
