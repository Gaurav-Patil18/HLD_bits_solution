// Problem: 45 - exams/m2014_q4i
module top_module (
    output out);
assign out=0;
endmodule
